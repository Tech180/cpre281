module Dflip_4bit(Q, D, EN, RST, CLK);
	input CLK, RST, EN;
	input [3:0] D;
	
	output [3:0] Q;

	wire [3:0] W1;
endmodule
